library verilog;
use verilog.vl_types.all;
entity CORDIC_vlg_vec_tst is
end CORDIC_vlg_vec_tst;

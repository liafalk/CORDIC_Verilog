// megafunction wizard: %Shift register (RAM-based)%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTSHIFT_TAPS 

// ============================================================
// File Name: shiftreg.v
// Megafunction Name(s):
// 			ALTSHIFT_TAPS
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 13.1.0 Build 162 10/23/2013 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2013 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module shiftreg (
	clock,
	shiftin,
	shiftout,
	taps);

	input	  clock;
	input	[31:0]  shiftin;
	output	[31:0]  shiftout;
	output	[63:0]  taps;

	wire [31:0] sub_wire0;
	wire [63:0] sub_wire1;
	wire [31:0] shiftout = sub_wire0[31:0];
	wire [63:0] taps = sub_wire1[63:0];

	altshift_taps	ALTSHIFT_TAPS_component (
				.clock (clock),
				.shiftin (shiftin),
				.shiftout (sub_wire0),
				.taps (sub_wire1)
				// synopsys translate_off
				,
				.aclr (),
				.clken ()
				// synopsys translate_on
				);
	defparam
		ALTSHIFT_TAPS_component.intended_device_family = "Cyclone III",
		ALTSHIFT_TAPS_component.lpm_hint = "RAM_BLOCK_TYPE=M9K",
		ALTSHIFT_TAPS_component.lpm_type = "altshift_taps",
		ALTSHIFT_TAPS_component.number_of_taps = 2,
		ALTSHIFT_TAPS_component.tap_distance = 6,
		ALTSHIFT_TAPS_component.width = 32;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ACLR NUMERIC "0"
// Retrieval info: PRIVATE: CLKEN NUMERIC "0"
// Retrieval info: PRIVATE: GROUP_TAPS NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
// Retrieval info: PRIVATE: NUMBER_OF_TAPS NUMERIC "2"
// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "1"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: TAP_DISTANCE NUMERIC "6"
// Retrieval info: PRIVATE: WIDTH NUMERIC "32"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
// Retrieval info: CONSTANT: LPM_HINT STRING "RAM_BLOCK_TYPE=M9K"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altshift_taps"
// Retrieval info: CONSTANT: NUMBER_OF_TAPS NUMERIC "2"
// Retrieval info: CONSTANT: TAP_DISTANCE NUMERIC "6"
// Retrieval info: CONSTANT: WIDTH NUMERIC "32"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: USED_PORT: shiftin 0 0 32 0 INPUT NODEFVAL "shiftin[31..0]"
// Retrieval info: USED_PORT: shiftout 0 0 32 0 OUTPUT NODEFVAL "shiftout[31..0]"
// Retrieval info: USED_PORT: taps 0 0 64 0 OUTPUT NODEFVAL "taps[63..0]"
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @shiftin 0 0 32 0 shiftin 0 0 32 0
// Retrieval info: CONNECT: shiftout 0 0 32 0 @shiftout 0 0 32 0
// Retrieval info: CONNECT: taps 0 0 64 0 @taps 0 0 64 0
// Retrieval info: GEN_FILE: TYPE_NORMAL shiftreg.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL shiftreg.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL shiftreg.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL shiftreg.bsf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL shiftreg_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL shiftreg_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf

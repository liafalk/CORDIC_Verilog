module CORDIC(
	theta,
	result
);

input wire	[31:0] theta;

ROM1	b2v_inst(
	
	.address(inputzz)
	);


endmodule
